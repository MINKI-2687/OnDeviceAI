module hello ();

endmodule
